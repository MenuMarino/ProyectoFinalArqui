module jump_and(input Branch, input Zero, output jump_and_out);

assign jump_and_out = Branch&Zero;

endmodule
